string
tasks[1] = '{"gen_data/task_1"};
